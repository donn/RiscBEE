`timescale 1ns/1ns

module BarrelShifter(A, O, shamt, arith, right);
    input [31:0] A;
    input [4:0] shamt;
    input arith, right;
    output [31:0] O;
    
    wire lastbit;
    assign lastbit = arith ? A[31] : 1'b0;
    
    genvar i, j;
    wire [31:0] C [5:0];
    
    //Use javascript.
    Mux2 #(1) mux0_0(.A(A[0]), .B(A[31]), .sel(right), .O(C[0][0]));
    Mux2 #(1) mux0_1(.A(A[1]), .B(A[30]), .sel(right), .O(C[0][1]));
    Mux2 #(1) mux0_2(.A(A[2]), .B(A[29]), .sel(right), .O(C[0][2]));
    Mux2 #(1) mux0_3(.A(A[3]), .B(A[28]), .sel(right), .O(C[0][3]));
    Mux2 #(1) mux0_4(.A(A[4]), .B(A[27]), .sel(right), .O(C[0][4]));
    Mux2 #(1) mux0_5(.A(A[5]), .B(A[26]), .sel(right), .O(C[0][5]));
    Mux2 #(1) mux0_6(.A(A[6]), .B(A[25]), .sel(right), .O(C[0][6]));
    Mux2 #(1) mux0_7(.A(A[7]), .B(A[24]), .sel(right), .O(C[0][7]));
    Mux2 #(1) mux0_8(.A(A[8]), .B(A[23]), .sel(right), .O(C[0][8]));
    Mux2 #(1) mux0_9(.A(A[9]), .B(A[22]), .sel(right), .O(C[0][9]));
    Mux2 #(1) mux0_10(.A(A[10]), .B(A[21]), .sel(right), .O(C[0][10]));
    Mux2 #(1) mux0_11(.A(A[11]), .B(A[20]), .sel(right), .O(C[0][11]));
    Mux2 #(1) mux0_12(.A(A[12]), .B(A[19]), .sel(right), .O(C[0][12]));
    Mux2 #(1) mux0_13(.A(A[13]), .B(A[18]), .sel(right), .O(C[0][13]));
    Mux2 #(1) mux0_14(.A(A[14]), .B(A[17]), .sel(right), .O(C[0][14]));
    Mux2 #(1) mux0_15(.A(A[15]), .B(A[16]), .sel(right), .O(C[0][15]));
    Mux2 #(1) mux0_16(.A(A[16]), .B(A[15]), .sel(right), .O(C[0][16]));
    Mux2 #(1) mux0_17(.A(A[17]), .B(A[14]), .sel(right), .O(C[0][17]));
    Mux2 #(1) mux0_18(.A(A[18]), .B(A[13]), .sel(right), .O(C[0][18]));
    Mux2 #(1) mux0_19(.A(A[19]), .B(A[12]), .sel(right), .O(C[0][19]));
    Mux2 #(1) mux0_20(.A(A[20]), .B(A[11]), .sel(right), .O(C[0][20]));
    Mux2 #(1) mux0_21(.A(A[21]), .B(A[10]), .sel(right), .O(C[0][21]));
    Mux2 #(1) mux0_22(.A(A[22]), .B(A[9]), .sel(right), .O(C[0][22]));
    Mux2 #(1) mux0_23(.A(A[23]), .B(A[8]), .sel(right), .O(C[0][23]));
    Mux2 #(1) mux0_24(.A(A[24]), .B(A[7]), .sel(right), .O(C[0][24]));
    Mux2 #(1) mux0_25(.A(A[25]), .B(A[6]), .sel(right), .O(C[0][25]));
    Mux2 #(1) mux0_26(.A(A[26]), .B(A[5]), .sel(right), .O(C[0][26]));
    Mux2 #(1) mux0_27(.A(A[27]), .B(A[4]), .sel(right), .O(C[0][27]));
    Mux2 #(1) mux0_28(.A(A[28]), .B(A[3]), .sel(right), .O(C[0][28]));
    Mux2 #(1) mux0_29(.A(A[29]), .B(A[2]), .sel(right), .O(C[0][29]));
    Mux2 #(1) mux0_30(.A(A[30]), .B(A[1]), .sel(right), .O(C[0][30]));
    Mux2 #(1) mux0_31(.A(A[31]), .B(A[0]), .sel(right), .O(C[0][31]));
    Mux2 #(1) mux1_0(.A(C[0][0]), .B(lastbit), .sel(shamt[4]), .O(C[1][0]));
    Mux2 #(1) mux1_1(.A(C[0][1]), .B(lastbit), .sel(shamt[4]), .O(C[1][1]));
    Mux2 #(1) mux1_2(.A(C[0][2]), .B(lastbit), .sel(shamt[4]), .O(C[1][2]));
    Mux2 #(1) mux1_3(.A(C[0][3]), .B(lastbit), .sel(shamt[4]), .O(C[1][3]));
    Mux2 #(1) mux1_4(.A(C[0][4]), .B(lastbit), .sel(shamt[4]), .O(C[1][4]));
    Mux2 #(1) mux1_5(.A(C[0][5]), .B(C[0][0]), .sel(shamt[4]), .O(C[1][5]));
    Mux2 #(1) mux1_6(.A(C[0][6]), .B(C[0][1]), .sel(shamt[4]), .O(C[1][6]));
    Mux2 #(1) mux1_7(.A(C[0][7]), .B(C[0][2]), .sel(shamt[4]), .O(C[1][7]));
    Mux2 #(1) mux1_8(.A(C[0][8]), .B(C[0][3]), .sel(shamt[4]), .O(C[1][8]));
    Mux2 #(1) mux1_9(.A(C[0][9]), .B(C[0][4]), .sel(shamt[4]), .O(C[1][9]));
    Mux2 #(1) mux1_10(.A(C[0][10]), .B(C[0][5]), .sel(shamt[4]), .O(C[1][10]));
    Mux2 #(1) mux1_11(.A(C[0][11]), .B(C[0][6]), .sel(shamt[4]), .O(C[1][11]));
    Mux2 #(1) mux1_12(.A(C[0][12]), .B(C[0][7]), .sel(shamt[4]), .O(C[1][12]));
    Mux2 #(1) mux1_13(.A(C[0][13]), .B(C[0][8]), .sel(shamt[4]), .O(C[1][13]));
    Mux2 #(1) mux1_14(.A(C[0][14]), .B(C[0][9]), .sel(shamt[4]), .O(C[1][14]));
    Mux2 #(1) mux1_15(.A(C[0][15]), .B(C[0][10]), .sel(shamt[4]), .O(C[1][15]));
    Mux2 #(1) mux1_16(.A(C[0][16]), .B(C[0][11]), .sel(shamt[4]), .O(C[1][16]));
    Mux2 #(1) mux1_17(.A(C[0][17]), .B(C[0][12]), .sel(shamt[4]), .O(C[1][17]));
    Mux2 #(1) mux1_18(.A(C[0][18]), .B(C[0][13]), .sel(shamt[4]), .O(C[1][18]));
    Mux2 #(1) mux1_19(.A(C[0][19]), .B(C[0][14]), .sel(shamt[4]), .O(C[1][19]));
    Mux2 #(1) mux1_20(.A(C[0][20]), .B(C[0][15]), .sel(shamt[4]), .O(C[1][20]));
    Mux2 #(1) mux1_21(.A(C[0][21]), .B(C[0][16]), .sel(shamt[4]), .O(C[1][21]));
    Mux2 #(1) mux1_22(.A(C[0][22]), .B(C[0][17]), .sel(shamt[4]), .O(C[1][22]));
    Mux2 #(1) mux1_23(.A(C[0][23]), .B(C[0][18]), .sel(shamt[4]), .O(C[1][23]));
    Mux2 #(1) mux1_24(.A(C[0][24]), .B(C[0][19]), .sel(shamt[4]), .O(C[1][24]));
    Mux2 #(1) mux1_25(.A(C[0][25]), .B(C[0][20]), .sel(shamt[4]), .O(C[1][25]));
    Mux2 #(1) mux1_26(.A(C[0][26]), .B(C[0][21]), .sel(shamt[4]), .O(C[1][26]));
    Mux2 #(1) mux1_27(.A(C[0][27]), .B(C[0][22]), .sel(shamt[4]), .O(C[1][27]));
    Mux2 #(1) mux1_28(.A(C[0][28]), .B(C[0][23]), .sel(shamt[4]), .O(C[1][28]));
    Mux2 #(1) mux1_29(.A(C[0][29]), .B(C[0][24]), .sel(shamt[4]), .O(C[1][29]));
    Mux2 #(1) mux1_30(.A(C[0][30]), .B(C[0][25]), .sel(shamt[4]), .O(C[1][30]));
    Mux2 #(1) mux1_31(.A(C[0][31]), .B(C[0][26]), .sel(shamt[4]), .O(C[1][31]));
    Mux2 #(1) mux2_0(.A(C[1][0]), .B(lastbit), .sel(shamt[3]), .O(C[2][0]));
    Mux2 #(1) mux2_1(.A(C[1][1]), .B(lastbit), .sel(shamt[3]), .O(C[2][1]));
    Mux2 #(1) mux2_2(.A(C[1][2]), .B(lastbit), .sel(shamt[3]), .O(C[2][2]));
    Mux2 #(1) mux2_3(.A(C[1][3]), .B(lastbit), .sel(shamt[3]), .O(C[2][3]));
    Mux2 #(1) mux2_4(.A(C[1][4]), .B(C[1][0]), .sel(shamt[3]), .O(C[2][4]));
    Mux2 #(1) mux2_5(.A(C[1][5]), .B(C[1][1]), .sel(shamt[3]), .O(C[2][5]));
    Mux2 #(1) mux2_6(.A(C[1][6]), .B(C[1][2]), .sel(shamt[3]), .O(C[2][6]));
    Mux2 #(1) mux2_7(.A(C[1][7]), .B(C[1][3]), .sel(shamt[3]), .O(C[2][7]));
    Mux2 #(1) mux2_8(.A(C[1][8]), .B(C[1][4]), .sel(shamt[3]), .O(C[2][8]));
    Mux2 #(1) mux2_9(.A(C[1][9]), .B(C[1][5]), .sel(shamt[3]), .O(C[2][9]));
    Mux2 #(1) mux2_10(.A(C[1][10]), .B(C[1][6]), .sel(shamt[3]), .O(C[2][10]));
    Mux2 #(1) mux2_11(.A(C[1][11]), .B(C[1][7]), .sel(shamt[3]), .O(C[2][11]));
    Mux2 #(1) mux2_12(.A(C[1][12]), .B(C[1][8]), .sel(shamt[3]), .O(C[2][12]));
    Mux2 #(1) mux2_13(.A(C[1][13]), .B(C[1][9]), .sel(shamt[3]), .O(C[2][13]));
    Mux2 #(1) mux2_14(.A(C[1][14]), .B(C[1][10]), .sel(shamt[3]), .O(C[2][14]));
    Mux2 #(1) mux2_15(.A(C[1][15]), .B(C[1][11]), .sel(shamt[3]), .O(C[2][15]));
    Mux2 #(1) mux2_16(.A(C[1][16]), .B(C[1][12]), .sel(shamt[3]), .O(C[2][16]));
    Mux2 #(1) mux2_17(.A(C[1][17]), .B(C[1][13]), .sel(shamt[3]), .O(C[2][17]));
    Mux2 #(1) mux2_18(.A(C[1][18]), .B(C[1][14]), .sel(shamt[3]), .O(C[2][18]));
    Mux2 #(1) mux2_19(.A(C[1][19]), .B(C[1][15]), .sel(shamt[3]), .O(C[2][19]));
    Mux2 #(1) mux2_20(.A(C[1][20]), .B(C[1][16]), .sel(shamt[3]), .O(C[2][20]));
    Mux2 #(1) mux2_21(.A(C[1][21]), .B(C[1][17]), .sel(shamt[3]), .O(C[2][21]));
    Mux2 #(1) mux2_22(.A(C[1][22]), .B(C[1][18]), .sel(shamt[3]), .O(C[2][22]));
    Mux2 #(1) mux2_23(.A(C[1][23]), .B(C[1][19]), .sel(shamt[3]), .O(C[2][23]));
    Mux2 #(1) mux2_24(.A(C[1][24]), .B(C[1][20]), .sel(shamt[3]), .O(C[2][24]));
    Mux2 #(1) mux2_25(.A(C[1][25]), .B(C[1][21]), .sel(shamt[3]), .O(C[2][25]));
    Mux2 #(1) mux2_26(.A(C[1][26]), .B(C[1][22]), .sel(shamt[3]), .O(C[2][26]));
    Mux2 #(1) mux2_27(.A(C[1][27]), .B(C[1][23]), .sel(shamt[3]), .O(C[2][27]));
    Mux2 #(1) mux2_28(.A(C[1][28]), .B(C[1][24]), .sel(shamt[3]), .O(C[2][28]));
    Mux2 #(1) mux2_29(.A(C[1][29]), .B(C[1][25]), .sel(shamt[3]), .O(C[2][29]));
    Mux2 #(1) mux2_30(.A(C[1][30]), .B(C[1][26]), .sel(shamt[3]), .O(C[2][30]));
    Mux2 #(1) mux2_31(.A(C[1][31]), .B(C[1][27]), .sel(shamt[3]), .O(C[2][31]));
    Mux2 #(1) mux3_0(.A(C[2][0]), .B(lastbit), .sel(shamt[2]), .O(C[3][0]));
    Mux2 #(1) mux3_1(.A(C[2][1]), .B(lastbit), .sel(shamt[2]), .O(C[3][1]));
    Mux2 #(1) mux3_2(.A(C[2][2]), .B(lastbit), .sel(shamt[2]), .O(C[3][2]));
    Mux2 #(1) mux3_3(.A(C[2][3]), .B(C[2][0]), .sel(shamt[2]), .O(C[3][3]));
    Mux2 #(1) mux3_4(.A(C[2][4]), .B(C[2][1]), .sel(shamt[2]), .O(C[3][4]));
    Mux2 #(1) mux3_5(.A(C[2][5]), .B(C[2][2]), .sel(shamt[2]), .O(C[3][5]));
    Mux2 #(1) mux3_6(.A(C[2][6]), .B(C[2][3]), .sel(shamt[2]), .O(C[3][6]));
    Mux2 #(1) mux3_7(.A(C[2][7]), .B(C[2][4]), .sel(shamt[2]), .O(C[3][7]));
    Mux2 #(1) mux3_8(.A(C[2][8]), .B(C[2][5]), .sel(shamt[2]), .O(C[3][8]));
    Mux2 #(1) mux3_9(.A(C[2][9]), .B(C[2][6]), .sel(shamt[2]), .O(C[3][9]));
    Mux2 #(1) mux3_10(.A(C[2][10]), .B(C[2][7]), .sel(shamt[2]), .O(C[3][10]));
    Mux2 #(1) mux3_11(.A(C[2][11]), .B(C[2][8]), .sel(shamt[2]), .O(C[3][11]));
    Mux2 #(1) mux3_12(.A(C[2][12]), .B(C[2][9]), .sel(shamt[2]), .O(C[3][12]));
    Mux2 #(1) mux3_13(.A(C[2][13]), .B(C[2][10]), .sel(shamt[2]), .O(C[3][13]));
    Mux2 #(1) mux3_14(.A(C[2][14]), .B(C[2][11]), .sel(shamt[2]), .O(C[3][14]));
    Mux2 #(1) mux3_15(.A(C[2][15]), .B(C[2][12]), .sel(shamt[2]), .O(C[3][15]));
    Mux2 #(1) mux3_16(.A(C[2][16]), .B(C[2][13]), .sel(shamt[2]), .O(C[3][16]));
    Mux2 #(1) mux3_17(.A(C[2][17]), .B(C[2][14]), .sel(shamt[2]), .O(C[3][17]));
    Mux2 #(1) mux3_18(.A(C[2][18]), .B(C[2][15]), .sel(shamt[2]), .O(C[3][18]));
    Mux2 #(1) mux3_19(.A(C[2][19]), .B(C[2][16]), .sel(shamt[2]), .O(C[3][19]));
    Mux2 #(1) mux3_20(.A(C[2][20]), .B(C[2][17]), .sel(shamt[2]), .O(C[3][20]));
    Mux2 #(1) mux3_21(.A(C[2][21]), .B(C[2][18]), .sel(shamt[2]), .O(C[3][21]));
    Mux2 #(1) mux3_22(.A(C[2][22]), .B(C[2][19]), .sel(shamt[2]), .O(C[3][22]));
    Mux2 #(1) mux3_23(.A(C[2][23]), .B(C[2][20]), .sel(shamt[2]), .O(C[3][23]));
    Mux2 #(1) mux3_24(.A(C[2][24]), .B(C[2][21]), .sel(shamt[2]), .O(C[3][24]));
    Mux2 #(1) mux3_25(.A(C[2][25]), .B(C[2][22]), .sel(shamt[2]), .O(C[3][25]));
    Mux2 #(1) mux3_26(.A(C[2][26]), .B(C[2][23]), .sel(shamt[2]), .O(C[3][26]));
    Mux2 #(1) mux3_27(.A(C[2][27]), .B(C[2][24]), .sel(shamt[2]), .O(C[3][27]));
    Mux2 #(1) mux3_28(.A(C[2][28]), .B(C[2][25]), .sel(shamt[2]), .O(C[3][28]));
    Mux2 #(1) mux3_29(.A(C[2][29]), .B(C[2][26]), .sel(shamt[2]), .O(C[3][29]));
    Mux2 #(1) mux3_30(.A(C[2][30]), .B(C[2][27]), .sel(shamt[2]), .O(C[3][30]));
    Mux2 #(1) mux3_31(.A(C[2][31]), .B(C[2][28]), .sel(shamt[2]), .O(C[3][31]));
    Mux2 #(1) mux4_0(.A(C[3][0]), .B(lastbit), .sel(shamt[1]), .O(C[4][0]));
    Mux2 #(1) mux4_1(.A(C[3][1]), .B(lastbit), .sel(shamt[1]), .O(C[4][1]));
    Mux2 #(1) mux4_2(.A(C[3][2]), .B(C[3][0]), .sel(shamt[1]), .O(C[4][2]));
    Mux2 #(1) mux4_3(.A(C[3][3]), .B(C[3][1]), .sel(shamt[1]), .O(C[4][3]));
    Mux2 #(1) mux4_4(.A(C[3][4]), .B(C[3][2]), .sel(shamt[1]), .O(C[4][4]));
    Mux2 #(1) mux4_5(.A(C[3][5]), .B(C[3][3]), .sel(shamt[1]), .O(C[4][5]));
    Mux2 #(1) mux4_6(.A(C[3][6]), .B(C[3][4]), .sel(shamt[1]), .O(C[4][6]));
    Mux2 #(1) mux4_7(.A(C[3][7]), .B(C[3][5]), .sel(shamt[1]), .O(C[4][7]));
    Mux2 #(1) mux4_8(.A(C[3][8]), .B(C[3][6]), .sel(shamt[1]), .O(C[4][8]));
    Mux2 #(1) mux4_9(.A(C[3][9]), .B(C[3][7]), .sel(shamt[1]), .O(C[4][9]));
    Mux2 #(1) mux4_10(.A(C[3][10]), .B(C[3][8]), .sel(shamt[1]), .O(C[4][10]));
    Mux2 #(1) mux4_11(.A(C[3][11]), .B(C[3][9]), .sel(shamt[1]), .O(C[4][11]));
    Mux2 #(1) mux4_12(.A(C[3][12]), .B(C[3][10]), .sel(shamt[1]), .O(C[4][12]));
    Mux2 #(1) mux4_13(.A(C[3][13]), .B(C[3][11]), .sel(shamt[1]), .O(C[4][13]));
    Mux2 #(1) mux4_14(.A(C[3][14]), .B(C[3][12]), .sel(shamt[1]), .O(C[4][14]));
    Mux2 #(1) mux4_15(.A(C[3][15]), .B(C[3][13]), .sel(shamt[1]), .O(C[4][15]));
    Mux2 #(1) mux4_16(.A(C[3][16]), .B(C[3][14]), .sel(shamt[1]), .O(C[4][16]));
    Mux2 #(1) mux4_17(.A(C[3][17]), .B(C[3][15]), .sel(shamt[1]), .O(C[4][17]));
    Mux2 #(1) mux4_18(.A(C[3][18]), .B(C[3][16]), .sel(shamt[1]), .O(C[4][18]));
    Mux2 #(1) mux4_19(.A(C[3][19]), .B(C[3][17]), .sel(shamt[1]), .O(C[4][19]));
    Mux2 #(1) mux4_20(.A(C[3][20]), .B(C[3][18]), .sel(shamt[1]), .O(C[4][20]));
    Mux2 #(1) mux4_21(.A(C[3][21]), .B(C[3][19]), .sel(shamt[1]), .O(C[4][21]));
    Mux2 #(1) mux4_22(.A(C[3][22]), .B(C[3][20]), .sel(shamt[1]), .O(C[4][22]));
    Mux2 #(1) mux4_23(.A(C[3][23]), .B(C[3][21]), .sel(shamt[1]), .O(C[4][23]));
    Mux2 #(1) mux4_24(.A(C[3][24]), .B(C[3][22]), .sel(shamt[1]), .O(C[4][24]));
    Mux2 #(1) mux4_25(.A(C[3][25]), .B(C[3][23]), .sel(shamt[1]), .O(C[4][25]));
    Mux2 #(1) mux4_26(.A(C[3][26]), .B(C[3][24]), .sel(shamt[1]), .O(C[4][26]));
    Mux2 #(1) mux4_27(.A(C[3][27]), .B(C[3][25]), .sel(shamt[1]), .O(C[4][27]));
    Mux2 #(1) mux4_28(.A(C[3][28]), .B(C[3][26]), .sel(shamt[1]), .O(C[4][28]));
    Mux2 #(1) mux4_29(.A(C[3][29]), .B(C[3][27]), .sel(shamt[1]), .O(C[4][29]));
    Mux2 #(1) mux4_30(.A(C[3][30]), .B(C[3][28]), .sel(shamt[1]), .O(C[4][30]));
    Mux2 #(1) mux4_31(.A(C[3][31]), .B(C[3][29]), .sel(shamt[1]), .O(C[4][31]));
    Mux2 #(1) mux5_0(.A(C[4][0]), .B(lastbit), .sel(shamt[0]), .O(C[5][0]));
    Mux2 #(1) mux5_1(.A(C[4][1]), .B(C[4][0]), .sel(shamt[0]), .O(C[5][1]));
    Mux2 #(1) mux5_2(.A(C[4][2]), .B(C[4][1]), .sel(shamt[0]), .O(C[5][2]));
    Mux2 #(1) mux5_3(.A(C[4][3]), .B(C[4][2]), .sel(shamt[0]), .O(C[5][3]));
    Mux2 #(1) mux5_4(.A(C[4][4]), .B(C[4][3]), .sel(shamt[0]), .O(C[5][4]));
    Mux2 #(1) mux5_5(.A(C[4][5]), .B(C[4][4]), .sel(shamt[0]), .O(C[5][5]));
    Mux2 #(1) mux5_6(.A(C[4][6]), .B(C[4][5]), .sel(shamt[0]), .O(C[5][6]));
    Mux2 #(1) mux5_7(.A(C[4][7]), .B(C[4][6]), .sel(shamt[0]), .O(C[5][7]));
    Mux2 #(1) mux5_8(.A(C[4][8]), .B(C[4][7]), .sel(shamt[0]), .O(C[5][8]));
    Mux2 #(1) mux5_9(.A(C[4][9]), .B(C[4][8]), .sel(shamt[0]), .O(C[5][9]));
    Mux2 #(1) mux5_10(.A(C[4][10]), .B(C[4][9]), .sel(shamt[0]), .O(C[5][10]));
    Mux2 #(1) mux5_11(.A(C[4][11]), .B(C[4][10]), .sel(shamt[0]), .O(C[5][11]));
    Mux2 #(1) mux5_12(.A(C[4][12]), .B(C[4][11]), .sel(shamt[0]), .O(C[5][12]));
    Mux2 #(1) mux5_13(.A(C[4][13]), .B(C[4][12]), .sel(shamt[0]), .O(C[5][13]));
    Mux2 #(1) mux5_14(.A(C[4][14]), .B(C[4][13]), .sel(shamt[0]), .O(C[5][14]));
    Mux2 #(1) mux5_15(.A(C[4][15]), .B(C[4][14]), .sel(shamt[0]), .O(C[5][15]));
    Mux2 #(1) mux5_16(.A(C[4][16]), .B(C[4][15]), .sel(shamt[0]), .O(C[5][16]));
    Mux2 #(1) mux5_17(.A(C[4][17]), .B(C[4][16]), .sel(shamt[0]), .O(C[5][17]));
    Mux2 #(1) mux5_18(.A(C[4][18]), .B(C[4][17]), .sel(shamt[0]), .O(C[5][18]));
    Mux2 #(1) mux5_19(.A(C[4][19]), .B(C[4][18]), .sel(shamt[0]), .O(C[5][19]));
    Mux2 #(1) mux5_20(.A(C[4][20]), .B(C[4][19]), .sel(shamt[0]), .O(C[5][20]));
    Mux2 #(1) mux5_21(.A(C[4][21]), .B(C[4][20]), .sel(shamt[0]), .O(C[5][21]));
    Mux2 #(1) mux5_22(.A(C[4][22]), .B(C[4][21]), .sel(shamt[0]), .O(C[5][22]));
    Mux2 #(1) mux5_23(.A(C[4][23]), .B(C[4][22]), .sel(shamt[0]), .O(C[5][23]));
    Mux2 #(1) mux5_24(.A(C[4][24]), .B(C[4][23]), .sel(shamt[0]), .O(C[5][24]));
    Mux2 #(1) mux5_25(.A(C[4][25]), .B(C[4][24]), .sel(shamt[0]), .O(C[5][25]));
    Mux2 #(1) mux5_26(.A(C[4][26]), .B(C[4][25]), .sel(shamt[0]), .O(C[5][26]));
    Mux2 #(1) mux5_27(.A(C[4][27]), .B(C[4][26]), .sel(shamt[0]), .O(C[5][27]));
    Mux2 #(1) mux5_28(.A(C[4][28]), .B(C[4][27]), .sel(shamt[0]), .O(C[5][28]));
    Mux2 #(1) mux5_29(.A(C[4][29]), .B(C[4][28]), .sel(shamt[0]), .O(C[5][29]));
    Mux2 #(1) mux5_30(.A(C[4][30]), .B(C[4][29]), .sel(shamt[0]), .O(C[5][30]));
    Mux2 #(1) mux5_31(.A(C[4][31]), .B(C[4][30]), .sel(shamt[0]), .O(C[5][31]));
    Mux2 #(1) mux6_0(.A(C[5][0]), .B(C[5][31]), .sel(right),   .O(O[0]));
    Mux2 #(1) mux6_1(.A(C[5][1]), .B(C[5][30]), .sel(right),   .O(O[1]));
    Mux2 #(1) mux6_2(.A(C[5][2]), .B(C[5][29]), .sel(right),   .O(O[2]));
    Mux2 #(1) mux6_3(.A(C[5][3]), .B(C[5][28]), .sel(right),   .O(O[3]));
    Mux2 #(1) mux6_4(.A(C[5][4]), .B(C[5][27]), .sel(right),   .O(O[4]));
    Mux2 #(1) mux6_5(.A(C[5][5]), .B(C[5][26]), .sel(right),   .O(O[5]));
    Mux2 #(1) mux6_6(.A(C[5][6]), .B(C[5][25]), .sel(right),   .O(O[6]));
    Mux2 #(1) mux6_7(.A(C[5][7]), .B(C[5][24]), .sel(right),   .O(O[7]));
    Mux2 #(1) mux6_8(.A(C[5][8]), .B(C[5][23]), .sel(right),   .O(O[8]));
    Mux2 #(1) mux6_9(.A(C[5][9]), .B(C[5][22]), .sel(right),   .O(O[9]));
    Mux2 #(1) mux6_10(.A(C[5][10]), .B(C[5][21]), .sel(right),   .O(O[10]));
    Mux2 #(1) mux6_11(.A(C[5][11]), .B(C[5][20]), .sel(right),   .O(O[11]));
    Mux2 #(1) mux6_12(.A(C[5][12]), .B(C[5][19]), .sel(right),   .O(O[12]));
    Mux2 #(1) mux6_13(.A(C[5][13]), .B(C[5][18]), .sel(right),   .O(O[13]));
    Mux2 #(1) mux6_14(.A(C[5][14]), .B(C[5][17]), .sel(right),   .O(O[14]));
    Mux2 #(1) mux6_15(.A(C[5][15]), .B(C[5][16]), .sel(right),   .O(O[15]));
    Mux2 #(1) mux6_16(.A(C[5][16]), .B(C[5][15]), .sel(right),   .O(O[16]));
    Mux2 #(1) mux6_17(.A(C[5][17]), .B(C[5][14]), .sel(right),   .O(O[17]));
    Mux2 #(1) mux6_18(.A(C[5][18]), .B(C[5][13]), .sel(right),   .O(O[18]));
    Mux2 #(1) mux6_19(.A(C[5][19]), .B(C[5][12]), .sel(right),   .O(O[19]));
    Mux2 #(1) mux6_20(.A(C[5][20]), .B(C[5][11]), .sel(right),   .O(O[20]));
    Mux2 #(1) mux6_21(.A(C[5][21]), .B(C[5][10]), .sel(right),   .O(O[21]));
    Mux2 #(1) mux6_22(.A(C[5][22]), .B(C[5][9]), .sel(right),   .O(O[22]));
    Mux2 #(1) mux6_23(.A(C[5][23]), .B(C[5][8]), .sel(right),   .O(O[23]));
    Mux2 #(1) mux6_24(.A(C[5][24]), .B(C[5][7]), .sel(right),   .O(O[24]));
    Mux2 #(1) mux6_25(.A(C[5][25]), .B(C[5][6]), .sel(right),   .O(O[25]));
    Mux2 #(1) mux6_26(.A(C[5][26]), .B(C[5][5]), .sel(right),   .O(O[26]));
    Mux2 #(1) mux6_27(.A(C[5][27]), .B(C[5][4]), .sel(right),   .O(O[27]));
    Mux2 #(1) mux6_28(.A(C[5][28]), .B(C[5][3]), .sel(right),   .O(O[28]));
    Mux2 #(1) mux6_29(.A(C[5][29]), .B(C[5][2]), .sel(right),   .O(O[29]));
    Mux2 #(1) mux6_30(.A(C[5][30]), .B(C[5][1]), .sel(right),   .O(O[30]));
    Mux2 #(1) mux6_31(.A(C[5][31]), .B(C[5][0]), .sel(right),   .O(O[31]));
    
endmodule 